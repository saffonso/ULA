library verilog;
use verilog.vl_types.all;
entity soma4bits_vlg_vec_tst is
end soma4bits_vlg_vec_tst;
