library verilog;
use verilog.vl_types.all;
entity soma4bits_vlg_check_tst is
    port(
        carry           : in     vl_logic_vector(1 downto 0);
        s               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end soma4bits_vlg_check_tst;
